LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE_232.ALL;
ENTITY CONTER IS 
	PORT (R : IN STD_LOGIC;
			E : IN STD_LOGIC;
			D : IN STD_LOGIC;
			Q : BUFFER STD_LOGIC;
			LDN : STD_LOGIC;
			RSTN : IN STD_LOGIC;
			UP_DNN : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			C : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE FUNC OF CONTER IS 
SIGNAL A0, A1, A2, A3, A4, A5, A6 : STD_LOGIC;
BEGIN 
U0 : XOR_2 PORT MAP (E, Q, A0);
M0 : MUX_2_1 PORT MAP (D, A0, LDN, A1);
M1 : MUX_2_1 PORT MAP (R, A1, RSTN, A2);
M2 : MUX_2_1 PORT MAP (A3, A4, UP_DNN, A5);
U1 : AND_2 PORT MAP (E, A5, C);
F0 : D_FF PORT MAP (A2, CLK, '1', '1', A3, A4);
q <= A3;
END FUNC;