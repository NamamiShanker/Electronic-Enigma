LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE_232.ALL;

ENTITY ELECTRONIC_ENIGMA_PRO IS
	PORT (I  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			D0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			D1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			D2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			LDNI : IN  STD_LOGIC;
			LDN  : IN STD_LOGIC;
			O   : INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			Q0  : INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			Q1  : INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			Q2  : INOUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			CLK : IN STD_LOGIC);
END ENTITY;

ARCHITECTURE FUNCTIONALITY OF ELECTRONIC_ENIGMA_PRO IS 
	
	SIGNAL Z0, Z1, Z2, Z3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL A0, A1, A2, A3, A4, A5: STD_LOGIC;
	BEGIN
	
		A0 <= I(0) OR I(1) OR I(2) OR I(3) OR I (4);
		A1 <= LDNI OR A0;
		C0 : COUNTER PORT MAP ("00000", D0, Q0, '1', LDN, '0', A1);
		A2 <= Q0(0) AND Q0(3) AND Q0(4);
		A3 <= LDNI OR A2;
		C1 : COUNTER PORT MAP ("00000", D1, Q1, '1', LDN, '0', A3);
		A4 <= Q1(0) AND Q1(3) AND Q1(4);
		A5 <= LDNI OR A4;
		C2 : COUNTER PORT MAP ("00000", D2, Q2, '1', LDN, '0', A5);

		M0 : MATCHER_1 PORT MAP (I, Z0);
		AR0: AR_CONV PORT MAP (Z0, Q0, Q1, CLK, Z1);
		M1 : MATCHER_2 PORT MAP (Z1, Z2);
		AR1: AR_CONV PORT MAP (Z2, Q1, Q2, CLK, Z3);
		M2 : MATCHER_3 PORT MAP (Z3, O);
	
END FUNCTIONALITY;


			
			
	
			