LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY XOR_2 IS
	PORT  (I0 : IN STD_LOGIC;
				 I1 : IN STD_LOGIC;
				 O0 : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE FUNC OF XOR_2 IS
BEGIN 
O0 <= I0 XOR I1;
END ARCHITECTURE;
